//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This sequences randomizes the inst_mem transaction and sends it 
// to the UVM driver.
//
// This sequence constructs and randomizes a inst_mem_transaction.
// 
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
class inst_mem_random_sequence 
  extends inst_mem_sequence_base ;

  `uvm_object_utils( inst_mem_random_sequence )

  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end
  
  //*****************************************************************
  function new(string name = "");
    super.new(name);
  endfunction: new

  // ****************************************************************************
  // TASK : body()
  // This task is automatically executed when this sequence is started using the 
  // start(sequencerHandle) task.
  //
  task body();
  
      // Construct the transaction
      req=inst_mem_transaction::type_id::create("req");
      start_item(req);
      // Randomize the transaction
      if(!req.randomize()) `uvm_fatal("SEQ", "inst_mem_random_sequence::body()-inst_mem_transaction randomization failed")
      // Send the transaction to the inst_mem_driver_bfm via the sequencer and inst_mem_driver.
      finish_item(req);
      `uvm_info("SEQ", {"Response:",req.convert2string()},UVM_MEDIUM)

  endtask

endclass: inst_mem_random_sequence

// pragma uvmf custom external begin
// pragma uvmf custom external end

