//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef enum bit [1:0] { CONTROL = 2'b00, DECODE = 2'b01, WRITEBACK = 2'b10, MEMORY = 2'b11 } block_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

