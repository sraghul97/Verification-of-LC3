//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef logic [15:0] vsr1_t;
typedef logic [15:0] vsr2_t;
typedef logic [2:0] psr_t;
typedef logic enable_writeback_out_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

